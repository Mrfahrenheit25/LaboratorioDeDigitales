03C28293800012B7
01C2A02300000E13
03828293800012B7
01C2802305500E13
4083031380001337
FFF38393000103B7
8000133700732023
000053B740430313
00010EB755538393
00400F93FFFE8E93
FFFF8F93020F8663
FFFF0F1300100F37
01D3C3B300732023
01DE4E3301C2A023
FFFF0F13FE0F00E3
800012B7FF9FF06F
00000E1303C28293
800012B701C2A023
00000E1303828293
8000133701C28023
0000039340430313
0000006F00732023
0000000000000000
